/*
    CS/ECE 552 Spring '20
    Homework #1, Problem 1

    1 input NOT
*/
module not1 (in1,out);
    input in1;
    output out;
    assign out = ~in1;
endmodule
